Komentar, naslov, ... prvo vrstico spice ignorira
    
    r_rs    3   6   r=5.4k
    r_rd    2   5   r=12.568k
    r_r1    3   4   r=37.5k
    r_r2    4   2   r=150.6k
    r_rsi   1   8   r=500
    r_rl    0   7   r=10k
    
    c_c1    8   4   c=100u
    c_c2    5   7   c=100u
    
    v_vin       1   0   dc=0    sin=(0,  0.012, 5k)
    v_vplus     3   0   dc=9
    v_vminus    2   0   dc=-9
    
    .model pmos1 pmos   level=1  vto=-0.5 kp=0.5m lambda=0
    
    
    m_m1    5   4   6   6   pmos1    w=15u    l=1u
    
    
    
    
    .control
        echo ########## Vaja 2 ##########
    
        echo .......... OP1 ..........
        
        op
           
            let idq=v(5,2) / 12568
            let vsdq=v(6,5)
            let vsgq=v(6,4)
            print idq vsdq vsgq
            
        
        echo .......... TRAN1 ..........
        
            tran  1u  5m
            let id=v(5,2) / 12568
            let vsd=v(6,5)
            let vsg=v(6,4)
            let vout=v(7)
            let vin=v(1)
            let vss=v(6)
            let vg=v(4)
            let vd=v(5)
            fourier 5k vout
            
            plot vss vg vd xlabel 'time' ylabel 'vs, vg, vd'
           
            let vin_pp=max(vin) - min(vin)
            let vout_pp=max(vout) - min(vout)
            let av=vout_pp/vin_pp
        
            print av
        
        
    .endc

    .end
