Naloga 2 
    * upornostni
    r_r1    1   2   r=37.5k
    r_r2    2   5   r=150.6k
    
    r_rs    1   3   r=5.432k
    r_rd    4   5   r=12.568k
    
    r_rsi	7	6	r=500
    r_rl	8	0	r=10k
    
    *kapacitivnosti
    c_c1	6	2	c=100u
    c_cs	3	0	c=100u
    c_c2	4	8	c=100u
    
    *napajalniki    
    v_vplus      1   0   dc=  9
    v_vminus     5   0   dc= -9
    v_in 		 7   0   dc=0    sin = (0, 0.0148, 5k)   
    
    *build our model
  	* m_imeTran d g s b (drain, gate, source, base) imeModela parametri
    * .model imeModela  tipElementa parametri(kp, vto, lambda,..)
    
    .model pmosTest pmos level=1 vto=-0.5 kp=0.5m
    m_ml    4   2   3   3   pmosTest    w=15u    l=1u
    
    .control
        destroy all
        
        echo _______________VAJA 2______________
        echo 
        
        *delovna tocka op -> poisce delovno tocko
        op
        
        echo _____________Naloga_2________________
        echo
        *nastavimo vektorje ki jih iscemo
        let idq  = v(1,3)/@r_rs[r]
        let vsdq = v(3,4)
        let vsgq = v(2,4)
        
        *izpis stevilk
        print idq vsdq vsgq 
        
        
        echo _____________Naloga_3________________
        echo "Sprememba kp poveca 10%"
        echo 
        
        idq_kp10posta = 5.027567e-04
        print idq_kp10posta 
        
        dIdq = idq_kp10posta/idq
        echo "Delta razlika Idq toka:"
        print dIdq
        
        echo _____________Naloga_4________________
        echo 
        
        tran 1u 5m
        	
        let id = v(1,3)/@r_rs[r]
		let vsd=v(3,4)
		let vsg=v(2,4)
		let vout=v(8)
		let vin=v(7)
		let vss=v(3)
		let vgg=v(2)
		let vdd=v(4)
		fourier 5k vout
		
		echo "plot"
        plot vss vgg vdd xlabel 'time' ylabel 'vs, vg, vd'
        
        
        *fourierova analiza
		echo _____________Naloga_5________________
        echo
        
			let vin_pp=max(vin)-min(vin)
			let vout_pp=max(vout)-min(vout)
			let av=vout_pp/vin_pp
			
			vs_pp=max(vss)-min(vss)
			vg_pp=max(vgg)-min(vgg)
			vd_pp=max(vdd)-min(vdd)
			
			plot vin vout
			print av vs_pp vg_pp vd_pp

          
      .endc
 .end

