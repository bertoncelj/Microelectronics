Vaja linel 2


vp 2 0 dc = 9
vm 5 0 dc = -9
vin 6 0 dc = 0	sin=(0, 0.01498, 5k)

r1 2 1 r=37.5k
r2 1 5 r=150.7k
rs 2 3 r=5.4k
rd 4 5 r=12.5k
rsi 6 7 r=500
rload 8 0 r=10k
c1 7 1 c=100u
c2 4 8 c=100u
*cs 3 0 c=100u

	*m_imeTran d g s b imeModela parametri
	*.model imeModela tipEl parametri(kp, vto, ...)

m1 4 1 3 3 modelp w=15u l=1u
	.model modelp pmos kp=0.5m vto=-0.5


.control
destroy all
    echo #### nal 2 ####

    
    echo ------OP1-------
	op
	let idq = v(2,3)/@rs[r]
	let vsdq = v(3,4)
	let vsgq = v(3,1)
	
	print idq vsdq vsgq 
	
	echo -----op2--------
    
    let @@modelp[kp] = 0.55m
 	op 
	let idq = v(2,3)/@rs[r]
	let vsdq = v(3,4)
	let vsgq = v(3,1)

	
    print idq vsdq vsgq
	
    let @@modelp[kp] = 0.5m
    op
	
	echo ------TRAN1------
	
        *tran dt            tstop
        *     časovni korak,konec
    tran 1u 3m
    fourier 5k v(8)
	
	plot v(1) v(4) v(3) xlabel 'time' ylabel 'vg, vd, vs' 
	*plot v(1) xlabel 'time' ylabel 'vgate[t]' 
	*plot v(4) xlabel 'time' ylabel 'vdrain[t]'
	*plot v(3) xlabel 'time' ylabel 'vsource[t]'
	plot v(8) v(6) xlabel 'time' ylabel 'vout[t], vin[t]'

	
	let vinPP = max(v(7))-min(v(7))
    let voutPP = max(v(8))-min(v(8))
    let avABS = voutPP/vinPP
    print avABS
    




.endc
 
.end
