Komentar,naslov... karkoli tukaj napisemo, spice ignorira, zadnja vrstica mora bita .end ce imamo ukaz .karkoli je to komanda simulatorju

* k-kilo, m-mili, meg-mega, u- mikro...
* masa je vedno vozlišče 0


*Opis vezja
* 1.crka: tip el. (r, c, l , m - mosfet, q- bjt,v,i...)
* sledi   : ime el.
* sledi   : vozl.
* sledi   : parametri

    rs 4    5   r = 4.38k
    rd 2    3   r = 8k
    
    *v_imeVira: n+ n- dc=xx acmag=xx sin=(offset,amplituda,frekvenca)
    vin 1   0   dc=0 sin= (0,1.3165834,1kHz)
    vdd 2   0   dc=5
    vss 0   5   dc=5

*   m_imeMosfeta d g s b imeModela parametri
* .model imeModela tipElementa parametri(kp,vto,lambda...)


    .model nmosTest nmos level=1 vto=1.4 kp=0.5m
    m1  3   1   4   4 nmosTest w=1u l=1u 

* komentar 
*ukazi:  echo, op, setplot, display, let, print, dc, tran
*Pri plotu lahko uporabimo vs -> Versus: Nariši vektor proti drugemu vektorju




.control
    destroy all
    echo ######## Vaja 1 ########
    
    
    ¸
    
    echo ............ OP1 .............
    *DelovnaTocka
    op
    
    *   print v(1) v(2) vin #branch i[v_vdd]
    * print all
    
    *Tok skozi tranzistor ID!
    *print -i(vdd) i(vss) v(2,3)/@rd[r]

    
    *spremenljivke (vektorji)
    
    let idq= -i(vdd)
    let vdsq=V(3,4)
    let vgsq = v(1,4)
    let vout=v(3)
    print idq vdsq vgsq vout
    
    echo ............ DC1 .............
    
    *dc analiza je serija op analiz
    *vector sweep zajema vrednosti, ki jih je dc spreminjal
    
    
    *dc param start stop korak
     dc @rs[r] 1k 10k 10
     
     *plot -i(vdd) xlabel 'RS[ohm]' ylabel 'IDQ[A]'
     
    echo ............ DC2 .............
    dc vin -10 10 0.01
    
    let id= -i(vdd)
    let vds=V(3,4)
    let vgs = v(1,4)
    let vout=v(3)
    
     *plot id vs vds xlabel 'vin[V]' ylabel 'Id[A]'
     *plot vout xlabel 'vin[V]' ylabel 'Vout[V]'
     
     echo ............ TRAN1 .............
     *tran dt tstop 
     tran 10u 5m
     
     let id= -i(vdd)
    let vds=V(3,4)
    let vgs = v(1,4)
    let vout=v(3)
     
     plot v(1) vout xlabel 'time' ylabel 'vin(t), vout(t)'
     
     * fourier popacenje
     * fourier f0 signal
     fourier 1k vout
     
     let vin_pp = max(v(1))-min(v(1))
     let vout_pp = max(v(3))-min(v(3))
     let av=vout_pp/vin_pp
     
     print av
    
.endc



.end
