 Komentar, naslov, opis vezja, ...
 
 * Komentar se začne z zvezdico in obsega celo vrstico
 
 * Opis vezja
 * Elementi:
 * 1. crka: Tip elementa (r, c, l, q, m, d, v, i, ...)
 * sledi: ime elementa
 * sledi: vozlisca
 * sledi: parametri
 
 r_rd           2   3   r=8k
 r_rs           4   5   r=4.37158k
 * Koncnice potenc 10: k-kilo, m-mili, meg-mega, u-mikro, g-giga, t-tera, n-nano
 * Brez enot

 * v_ime        n+  n-  dc=xxx sin=(offset, amplituda, frekvenca)   acmag=xxx
 v_vin          1   0   dc=0    sin=(0, 10, 1k)
 v_vdd          2   0   dc=5
 v_vss          5   0   dc=-5
 
 * Mosfet
 * m_ime        drain   gate   source   bulk    ime_modela  parametri
 m_m1           3       1      4        4       testmodel   w=2u l=1u
 
* model: .model ime_modela tip_elementa parametri (kp parameter je v ucbeniku kp')
 .model     testmodel   nmos    vto=1.4     kp=0.25m     lambda=0
* Kontrol blok, notri so ukazi
* Ukazi: echo (izpiše tekst v okno simulatorja)
*        cd (zamenja mapo)
*        op (analiza delovne tocke)
*        setplot
*        destroy (all ali posamezno)
*        display (pokaze kaj je SPICE izracunal v zadnji analizi)
*        i(ime vira) (dostop do toka skozi vir)
*        let (to je za delat s spremenljivkami)
*        dc (dc analiza)
*        plot ()
*        tran
*        fourier
*        max (maksimalna vrednost)
*        min (minimalna vrednost)




 .control
    destroy all
    echo ########################## START ###########################
    echo --------------------------__OP1__---------------------------
    op
    
    *IDQ: vRD/RD =v(2,3)/rd
    *print -i(v_vdd)     v(2,3)/@r_rd[r]   v_vss#branch
    
    let idq=-i(v_vdd)
    let vdsq=v(3,4)
    let vgsq=v(1,4)
    let vout=v(3)
    
    print idq vdsq vgsq vout
    
    echo --------------------------__DC1__---------------------------
    * dc parameter start stop korak
    dc @r_rs[r] 1k 10k 10
    
    let idq=-i(v_vdd)
    let vdsq=v(3,4)
    let vgsq=v(1,4)
    let vout=v(3)
    
    *plot idq xlabel 'Rs [Ohm]' ylabel 'IDQ [A]'
    *plot -i(v_vdd)
    
    echo --------------------------__DC1__---------------------------
    *dc @v_vin[dc] -10 10 1 ista stvar kot naslednja vrstiva
    dc v_vin -10 10 0.1
    
    let id=-i(v_vdd)
    let vds=v(3,4)
    let vgs=v(1,4)
    let vout=v(3)
    
    *plot id vs vds xlabel 'vin [V]' ylabel 'id [A]'
    *plot vout vs sweep xlabel 'vin [V]' ylabel 'vout [V]'
    
    echo --------------------------_TRAN1_---------------------------
    * tran dt tstop
    tran    10u 5m
    
    let id=-i(v_vdd)
    let vds=v(3,4)
    let vgs=v(1,4)
    let vout=v(3)
    let vin=v(1)
    
    plot vin vout xlabel 'time' ylabel 'r:vin, g:vout'
    
    * Analiza popačenja Fourierova analiza
    * fourier f0 signal
    fourier 1k vout
    
    let vin_pp=max(vin)-min(vin)
    let vout_pp=max(vout)-min(vout)
    let av_abs=vout_pp/vin_pp
    print av_absz
    
 .endc
 .end
 
 
 * Dostop do vaj od doma: lisa.fe.uni-lj.si/vaje    Uporabnik: vaje Geslo: vajenec
