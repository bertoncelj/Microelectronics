 Komentar, naslov, Vaja1
    

 r_r1   1   2  r=1k
 r_r2   3   0  r=2k
 c_c1   2   3  c=1u
 c_c2   3   0  c=0.1n
 *acmag rabmo za ac analizo
 v_vin  1   0   dc=0  sin=(1, 1, 1k) acmag=1

 

 
 .control
    destroy all
    
    echo #########
    *malosignalna izmenicna analiza => potrebuje vsaj en acmag vir, pol sinus zravn nima veze
    *ac tip_skale(lin, log) st_tock_na_dekado fstart fstop
    ac dec 10 1 100meg
   
   let av=v(3)/v(1)
   let av_db=db(av)
   let av_ph=ph(av)
   plot av_db xlabel 'f' ylabel 'Av[dB]'
   plot av_ph xlabel 'f' ylabel 'Ph'
 .endc
                 
 .end
