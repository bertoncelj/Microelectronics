vaja 4
 .include models.inc
 r_rsrc 0 2 r=10k
 r_r1   3 4 r=242k
 r_r2   3 6 r=395k
 r_re   5 6 r=10k
 *r_rl   7 0 r=20k
 

 c_c1   2 3 c=100u
 c_c2   5 7 c=100u
 
 v_vp   4 0 dc=5
 v_vn   6 0 dc=-5
* v_vsrc 1 0 dc=0    sin(0,1,5k)
 v_vmer1    3 8 dc=0
 v_vmer2    9 4 dc=0
 v_Vx 7 0 dc=0 sin(0,2,5k)

 
 

 Q_Q1 (9 8 5) BC238B
 
 
 
 
 
 
 
 
 .control
    
    destroy all
    
    echo ##################### Vaja 4 ############################
    
    
    echo --------------------------------transientna analiza----------------------------------
    
    tran 1u 0.5m
    
    let Ix=i(v_vx)
   
    
    let Vx_pp=max(v(7))-min(v(7))
    let Ix_pp=max(Ix)-min(Ix)

    let Rout=Vx_pp/Ix_pp

    print Rout
    
  

    
    
    .endc
    
.end
    
   