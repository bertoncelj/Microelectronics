Komentar, opis, naslov,...
 
 
*komentar se začne z zvezdico
 
*opis vezja 
*elementi:
*1. crka: tip elementa(r,c,l,q,n,d,v,i,...)
*   sledi: ime elementa
*   sledi: vozlišča
*   sledi: parametri

* ignorira velike in male črke
* koncnice potenc 10 (k-kilo, m-mili, meg-mega, u-mikro, g, t, n, f,...)
* brez enot
r_rd            2   3   r=8k
r_rs            4   5   r=4.4k

*najprej + potem - vozlišče, dc=xxx sin(offset, ampl, frekvenca), acmag=xxx
v_vin           1   0   dc=0           sin(0,0.5,1K)
v_vdd           2   0   dc=5
v_vss           5   0   dc=-5

*  mosfet tranzistor
*m_ime d g s b (drain gate source bulk) ime_modela parametri
m_m1            3  1   4   4   testmodel w=2u l=1u

*model: .model ime_modela tip_elementa parametri
 .model testmodel nmos vto=1.4 kp=0.25m lambda=0
 
 
 
 
 
*kontrol blok-ukazi
*ukazi: echo, op, setplot, destroy, display, print, let, dc, plot, tran, fourier, max, min

.control
    destroy all
    echo ####################    START    ##########################
 
    echo ------------------OP--------------------------------
    op
   *IDQ, vRD/RD=v(2,3)/rd
  * print -i(v_vdd)  v(2,3)/@r_rd[r] v_vss#branch
   
   let idq=-i(v_vdd) 
   let vdsq=v(3,4)
   let vgsq=v(1,4)
   let vout=v(3)
   print idq vdsq vgsq vout
   
   *enosmerna analiza
   echo -----------------------DC1------------------------------------
   *dc parameter start stop korak
   dc @r_rs[r] 1k 10k 10
   
   let idq=-i(v_vdd) 
   let vdsq=v(3,4)
   let vgsq=v(1,4)
   let vout=v(3)
   
  * plot idq xlabel 'RS[ohm]' ylabel 'IDQ [A]'
 
  echo -----------------------DC2------------------------------------
  *dc @v_vin[dc] -10 10 1
  dc v_vin -10 10 0.1
  let id=-i(v_vdd) 
   let vds=v(3,4)
   let vgs=v(1,4)
   let vout=v(3)
  
  
 * plot id vs vds xlabel 'vds[V]' ylabel 'id[A]'
 * plot vout xlabel 'vin[V]' ylabel 'vout[V]'
 
 
 echo -----------------------tran1-------------------------------
 *tran dt tstop

 tran 1u 5m
  let id=-i(v_vdd) 
   let vds=v(3,4)
   let vgs=v(1,4)
   let vout=v(3)
   let vin =v(1)
 
 plot vin vout  xlabel 'table' ylabel 'r:vin,g:vout'
 
 * fourier analiza popačenja
 * fourier f0 signal
 fourier 1k vout
 
 let vin_pp=max(vin)-min(vin)
  let vout_pp=max(vout)-min(vout)
 let av_abs=vout_pp/vin_pp
print av_abs
 
 
 
 
 
 
 
 
 
 
 
 
 
 
.endc
.end
