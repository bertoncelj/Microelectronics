Komentar, naslov,..... (1 vrstico SPICE ingnorira)
    *VSE Z MALO
    
    * Opis vezja
    * 1.crka: tip elementa (r, c, l, m -mosfet, q-bjt, v -napetostni vir, i-* tokovni vir)
    * sledi  : ime el.
    * sledi   : vozel
    *sledi      : parametri
    
    *faktorji multiplikacije
    * k-kilo, m-mili, meg -mega, u-mikro,...
    
    *masa je vedno vozlišče nic
    *ce rabis ket tok zmerit urens notri napajlnik
    *sweep je default scale-> nvm googli neki pomembenga
    
    *v_imevira za napetostne vire n+, n- 
    *parametri za napajalnik
        *dc=xx
        *acmag=xx sin= (offset, ampl, freq)
    
    r_rs    4   5   r=4.4k
    r_rd    2   3   r=8k
    
    v_in    1   0   dc=0    sin = (0, 1.3, 1k)    
    v_vdd   2   0   dc=5
    v_vss   5   0   dc=-5
            
    * m_imeTran d g s b (drain, gate, source, base) imeModela parametri
    * .model imeModela  tipElementa parametri(kp, vto, lambda,..)

    .model nmosTest nmos level=1 vto=1.4 kp=0.5m
    m_ml    3   1   4   4   nmosTest    w=1u    l=1u
    
    
    
    *Ukazi:
    *   echo: izpis + locimo med izpisi
    *   op: resi enacbo
    *   setplot: napises v spiceopus da ti da vn kakšne je opravil
    *   display: katere stevilke je spice zracunob
    *   let: isto kot display
    *   print: 
    *   let 
    *   dc
    *   destroy
    *   plot
    *   tran
    *   fourier
    *   max, min 
    
    .control
        echo Hello World
        echo /************** VAJA 1 ******************/
        *pobrisemo vse spremeljivke, prosti polnilnik
        destroy all
        
        
        
        
        
        *delovna tocka op -> poisce delovno tocko
        op
        
        *print v(1) v(2) v_in#beanch
        * print all
        
        * tok skozi tranzistor
        print -i(v_vdd) i(v_vss)    v(2,3)/@r_rd[r]
        
        *spremeljivke (vektorji)
        let idq=i(v_vss)
        let vdsq =v(3,4)
        let vgsq = v(1,4)
        let vout = v(3)
        print idq vdsq vgsq vout
        
        print idq, vdsq, vgsq
        
        echo ........DC ANALIZA............
        * enosmerna analiza
        * dc param start stop korak
        *tako spreminajmo en paramater z @
        dc @r_rs[r] 1k 10k 10
        
        *plot -i(v_vdd) xlabel 'RS[ohm]' ylabel 'IDQ [A]'
        
        echo .................DC 2...................
        *tukaj bi tudi mogli pisat @ ampak ne rabmo
        dc v_in -10 10 0.1
        
        let id= -i(v_vdd)
        let vds = v(3,4)
        let vgs = v(1,4)
        let vout = v(3)
        
        *vs pomeni neki proti neki ce hocs popravit default skalo
        *plot id vs vds xlabel 'vds[V]' ylabel 'id[A]'
        
        *plot vout xlabel 'vin[V]' ylabel 'vout[V]'
        
        *za 4 nalogo kliknes na grafu in pogledas odvod da dobis koificjen
        
         echo .................TRANZIANT ANALYSIS...................
         *  tran dt tstop -> najbolj osnovna verzija
         *     - dt je korak 
         *     - tstop koliko signaala zahtevamo
         tran 10u 5m 
         
         let id= -i(v_vdd)
         let vds = v(3,4)
         let vgs = v(1,4)
         let vout = v(3)
        
         plot v(1) vout xlabel 'time [s]' ylabel 'r:vin(t), g:vout(t)'
         
         *  fourier analiza za popacenje
         *  fourier f0 signal ->syntakse
         fourier 1k vout
         
         let vin_pp = max(v(1)) - min(v(1))
            let vout_pp = max(v(3)) - min(v(3))
         let av = vout_pp/vin_pp
         print av
         *manka av minus ker je v protifazi
    .endc
    
    .end
