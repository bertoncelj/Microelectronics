Ime

    .control
    
    .endc
    
.end
