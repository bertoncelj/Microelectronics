Emitorski sledilnik - izhodna upornost
.include models.inc

vin 1 0 dc = 0 
vp 6 0 dc = 5
vn  4 0 dc = -5
voutt 7 0 dc = 0 sin(0 1 5k)

r1 6 3 r=175k
r2 3 4 r=216k
re 4 5 r=6.415k

rsrc 1 2 r=10k

q1 6 3 5 BC238B

c1 2 3 c=100u
c2 5 7 c=100u


.control
tran 1u 3m
let ix = max(i(voutt)) - min(i(voutt))
let vx = max(v(7))-min(v(7))
let rout = vx/ix
print rout


.endc
.end
