.control
    destroy all
    echo ########### Vaja * ###########
    
    
    
    
    
    
    
    
    
    

.endc
.end  
