Komentar, naslov, opis,....

* komentar se zacne z


* Opis vezja
* elementi:
*   1.crka: tip el. (r, c, l, q, m, d, v, i, ...)
*   sledi:  ime el. 
*   sledi:  vozl. 
*   sledi:  parametri

* koncnice potenc 10: k-kilo, m-mili, meg-mega, u-mikro, g, t, n, p, f,
* brez enot

r_rd        2   3   r=8k
r_rs        4   5   r=4.4k

*v_ime      n+  n-  dc=xxx sin=(offset, ampl, ferkv)  acmag=xxx
v_vin       1   0   dc=0    sin=(0, 1.0, 1k)
v_vdd       2   0   dc=5
v_vss       5   0   dc=-5


*mosfet
* mime  drain gate source bulk  ime_modela parametri
m_m1        3   1   4   4   testmodel w=2u l=1u 

*model: .model ime_modela tip_el parametri
.model testmodel nmos vto=1.4 kp=0.25m lambda=0





* kontrol block - ukazi
* ukazi: echo, op, seplot, destroy, display, print, let, dc, plot, tran, fourier, max, min

.control
    destroy all

    echo ###################### START ################

    echo -------------------- OP1 --------------------
    op
    
    *IDQ: vRD/RD = v(2,3)/rd
    * print -i(v_vdd)  v(2,3)/@r_rd[r]  v_vss#branch
    
    let idq=-i(v_vdd)
    let vdsq=v(3,4)
    let vgsq=v(1,4)
    let vout=v(3)
    
    print idq vdsq vgsq vout
    
    
    * enosmerna analiza
    echo ------------------ DC1 -----------------
    * dc param start stop korak
    dc @r_rs[r] 1k 10k 10
    
    let id=-i(v_vdd)
    let vds=v(3,4)
    let vgs=v(1,4)
    let vout=v(3)

    *plot id  xlabel 'RS [ohm]' ylabel 'IDQ [A]'
    
    
    echo ------------------ DC2-----------------
    *dc @v_vin[dc] -10 10 1
    dc v_vin -10 10 0.1
    
    let id=-i(v_vdd)
    let vds=v(3,4)
    let vgs=v(1,4)
    let vout=v(3)

    
    *plot id vs vds xlabel 'vds[V]' ylabel 'id[A]' 
    *plot vout xlabel 'vin[V]' ylabel 'vout[V]' 
    
    
    echo ------------------ TRAN1 -----------------
    * tran dt tstop
    tran 1u 5m

    
    let id=-i(v_vdd)
    let vds=v(3,4)
    let vgs=v(1,4)
    let vout=v(3)
    let vin=v(1)
    
    plot vin vout xlabel 'time' ylabel 'r:vin, g:vout'
    
    
    *fourier  - analiza popacenja
    * fourier f0 signal
    fourier 1k vout
    
    let vin_pp=max(vin)-min(vin)
    let vout_pp=max(vout)-min(vout)
    let av_abs=vout_pp/vin_pp
    print av_abs
    
.endc
.end

