Komentar, naslov, opis... spice opus to vedno ignorira

* komentar se zacne z zvezdico - cela vrstica ignorirana

* spice ni case-sensitive... M=m

* opis vezja - pred kontrol blokom - elementi vezja - spice dela z vozlisci 
* elementi:
*   1. crka = tip el. (r, c, l, q, m, d, v, i, ...)
*   sledi: ime el. 
*   sledi: vozlisca
*   sledi: parametri
*   spice prepoznava koncince potenc 10: k-kilo, m-mili, meg-mega, u-mikro
*                                        g-giga, t-tera, n-nano itd...
* BREZ ENOT, samo koncnice!

r_rd    2   3   r=8k
r_rs    4   5   r=4.4k

*v_ime +vozlisce -vozlisce dc=xxx sin=(offset, ampl, frekv) acmag=xxx 
v_vin   1   0   dc=0 sin=(0, 1.0, 1k)
v_vdd   2   0   dc=5
v_vss   5   0   dc=-5

* mosfet
*m_ime d (drain) g (gate) s (source) b (bulk - substrat) ime_mod parametri
*m_ime d g s b 

m_m1    3   1   4   4   testmodel  w=2u l=1u  

*model: .model ime_modela tip_elementa parametri

.model  testmodel   nmos    vto=1.4     kp=0.25m lambda=0

* default w/l=1
*kp = k' v nasi literaturi



* kontrol blok - tuki not bojo ukaz ki jih izvaja simulator
* ukazi: echo (izpis teksta v simulator), op (analiza delovne tocke)
*        setplot(poglej vse analize za nazaj), destroy all (izbrisi vse)
*        display (rezultati anazlize - potenciali, #branch -> tokovi virov
*        print (stevilska vrednost spremenljivk), let (spremenljivka)
*        dc (dc analiza), plot, tran - tranzienta analiza, fourier, max,
*        min

* CE IMAMO DIODO DODAMO NAPETOSTI VIR ZAPOREDNO Z DC=0 in SPICE zracuna tok

.control

    destroy all

    echo ### START ###
    
    echo ----- OP1 -----
    op
    *IDQ - vRD/RD = v(2,3)/RD -- [r] <- paramter r (upornost)
    *print -i(v_vdd) v(2,3)/@r_rd[r] v_vss#branch NI PREGLEDNO
    
    *let - spremenljivk
    
    let idq=v_vss#branch 
    let vdsq=v(3,4)
    let vgsq=v(1,4)
    let vout = v(3)
    
    print idq vdsq vgsq vout
    
    echo ------------------- DC analiza 1 ------------------------
    * polgej enosmerne razmere za razlicne parametre
    * dc paramter_spremenljiv start stop korak
    
    dc @r_rs[r] 1k 10k 10
    
    let idq=v_vss#branch 
    let vdsq=v(3,4)
    let vgsq=v(1,4)
    let vout = v(3)
    
    *plot idq xlabel 'RS[ohm]' ylabel 'IDQ [A]'
    
    echo ------------------- DC analiza 2 ------------------------
    
    *spreminjamo v_vin (dc) po 1 volt med -10 do 10
    
    *dc @v_vin[dc] -10 10 1 --> isto kot psondje ker ze ima dc parameter
    
    
    dc v_vin -10 10 0.1
    
    let id=v_vss#branch 
    let vds=v(3,4)
    let vgs=v(1,4)
    let vout = v(3)
    let vin = (v1)
    
    *plot id vs vds xlabel 'vds[V]' ylabel 'id[A]'
    
    *plot vout vs sweep xlabel 'vin[V]' ylabel 'vout[V]'
    
    echo ------------------- TRAN1 ------------------------
    * tran dt tstop
    
    tran 1u 5m
    
    let id=v_vss#branch 
    let vds=v(3,4)
    let vgs=v(1,4)
    let vout = v(3)
    let vin = v(1)
    
    plot vin vout xlabel 'time' ylabel 'r:vin, g:vout'
    
    * fourier - analiza popacenja
    * fourier f0 signal
    
    fourier 1k vout
    
    let vin_pp=max(vin)-min(vin)
    let vout_pp=max(vout)-min(vout)
    let av_abs=vout_pp/vin_pp
    print av_abs
    
    
.endc

.end
