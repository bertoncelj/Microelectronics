Vaja linel 3 


vp 4 0 dc = 5
vn 8 0 dc = -5
vin 1 0 dc = 0	sin=(0, 0.0, 5k)
vout 9 0        sin=(0, 0.2, 5k)

r1 3 4 r=40.484k
r2 2 3 r=31.628k
r3 8 2 r=54.4k
rs 7 8 r=5k
rd 4 5 r=5k

c1 1 2 c=100u
c2 3 0 c=100u
c3 7 0 c=100u
c4 5 9 c=100u

	*m_imeTran d g s b imeModela parametri
	*.model imeModela tipEl parametri(kp, vto, ...)

.model modeln nmos kp=0.5m vto=0.8 lambda=0.1m

m1 6 2 7 7 modeln w=2u l=1u
m2 5 3 6 6 modeln w=2u l=1u	
	

.control
destroy all
    
	
        tran 1u 5m
  
        
        let voutPP = max(v(9))-min(v(9))
        let ioutPP = max(i(vout))-min(i(vout))
        let rout = voutPP/ioutPP
        print rout
        
        

.endc
 
.end
