


vx 1 0 dc=0 sin=(0, 1, 1k)
r1 1 2 r=1k
r2 2 0 r=2k




.control
destroy all

*tf out vir


.endc
.end 
