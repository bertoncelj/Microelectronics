Uvod pri vaji  5: ac analiza

vin 1 0 dc= 0 sin = (1, 1, 1k), acmag= 1
*acmag rabimo pri ac analizi, vsaj en acmag vir!!
r1 1 2 r=1k
c1 2 3 c=1u
r2 3 0 r=2k
c2 3 0 c=0.1n

.control
destroy all

echo #####################################################

*malosignalna izmenična analiza 
* sintaksa: ac tip_skale st_tock fstart f stop ( dec - dekada, logaritemska skala, f start stop = začetna in končna frekvenca) 

ac dec 10 1 100meg

let av=v(3)/v(1)
let av_db = db(av)  
let av_ph = ph(av)  

* decibeli db
*ph kot faza

plot av_db xlabel 'f' ylabel 'av[dB]'
plot av_ph xlabel 'f' ylabel 'phase'




.endc
.end
