 Design Example 6.7
	r_rc	3	4	r=10k
	r_rb	2	3	r=100k
	
	r_re1	5	6	r=240
	r_re2	6	7	r=20k	

*napajniki
	
	v_vplus 	3	0	dc= 5
	v_vminus	7	0	dc=-5	
	v_vs		1	0	dc= 0	sin = (12m, 0.0148, 2k)

*kondez
	c_c1	1	2	c=100u
	c_c5	6	0	c=100u

  *includamo tranzistor
    .include models.inc
  
  * m_imeTran (c b e) imeModela parametri
    q_q1    4 2 5 5  T2N2222
    
    .control
    destroy all
           
    echo _________Example 6.7__________
    echo
    echo        
    echo .........Preverimo delovno tocko.........
       
    *naredi DC analizo
    op
            
    *nastavimo vektorje ki jih iscemo
    let icq   = v(3,4)/@r_rc[r]
    
            
    *izpisemo vektroje
     print icq
    
     
    echo 
    echo .........NALOGA_3................
     
    echo ----------------------Napetostno, Tokovno ojacanje-----------------------------
	
	tran 1u 5m
	
	*napetostno ojacanje
		let vout=v(4)
		let vin=v(1)

    	let vout_pp=max(vout)-min(vout)
		let vin_pp=max(vin)-min(vin)
	
		let Av = vout_pp/vin_pp
		
	*izpise ojacanje
	print  Av

    
    .endc
    
.end
