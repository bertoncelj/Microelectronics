Naslov vaje


.control


.endc


.end
