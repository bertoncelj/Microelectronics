 
  *****Labvaja3******


  *opis vezja
  *1.crka     :tip el. (r,c,l,m -mostfet, q-bjt, v,i,...)
  *sledi      : ime el.
  *sledi      : vozl.
  *sledi      :parametri
  
  
  *masa: vozlisce 0
  *k-kilo, m-mili, meg - mega, u-mikro,...
  
  
  rs     (7  8)   r=5k
  rd     (4  5)   r=5k
  r1     (4  3)   r=45.6k
  r2     (3  2)   r=35.63k
  r3     (2  8)   r=61.28k
  
  
  cl     (1  2)   c=100u
  c2     (0  3)   c=100u
  c3     (7  0)   c=100u
  c4     (5  10)   c=100u
  
  
  *v:imevira n+ n-  dc=xx acmag=xx  sin(offset, amplituda, frekvenca) 
  
  vin   (1  0)  dc=0   sin=( 0, 0, 0)
  vnn   (8  0)  dc=-5
  vpp   (4  0)  dc=5
  vgg   (10 0)  dc=0   sin=( 0, 0.04, 5k) 
  
  
  
  *m imeTranzistorja  d g  s c imeModela parametri
  * .model imeModela tipEl parametri(kp,vto, labda...)
  
  
  .model nmosTest nmos level=1  vto=0.8 kp=1m lambda= 0.1m
  
  m1  (6  2  7  7)   nmosTest  w=1  l=1
  m2  (5  3  6  6)   nmosTest  w=1  l=1
  
  
  

 *komentar
 *ukazi: echo, op, setplot, display, print, let ,dc, destroy, plot, tran, fourier, max, min, sqrt
 
 

  .control
     destroy all
    echo  ################################Vaja 3##################################
     
     
     echo  .................................OP1.....................................
     *delovna tocka
     op
     
     * print v(1), print v(2), print all, print vdd#branch,...
     
     
     
     
     *spremenljivke (vektorji)
     
     let idq= v(4,5)/@rd[r]
     print idq
     
     let vds2q= v(5,6)
     let vds1q= v(6,7)
     let vgs2q= v(3,6)
     let vgs1q= v(2,7)
     let vg1=v(1)
     let vout=v(5)
     print  vds1q vds2q  vgs1q  vgs2q vout vg1
     
     
    
     
     
    
     
      echo .............. TRAN0.............
     *tran dt tstop
     
     tran 0.005u 1m
     
     let idq= v(4,5)/@rd[r]
   
     
     let vds2q= v(5,6)
     let vds1q= v(6,7)
     let vgs2q= v(3,6)
     let vgs1q= v(2,7)
     let vg1=v(1)
     let vout=v(5)
     
     
     
     *plot v(1) vss xlabel 'time' ylabel 'r:vin(t), g:vs(t)'
     *plot v(1) vg xlabel 'time' ylabel 'r:vin(t), g:vg(t)'
     *plot v(1) vd xlabel 'time' ylabel 'r:vin(t), g:vd(t)'
     
     *plot vout vs vin xlabel 'vin' ylabel 'r:vout'
     
    *plot v(1) vout vss vg vd  xlabel 'time' ylabel 'r:vin(t), g:vout(t), b:vs(t), g:vg(t), k:vd(t)'
    
      
      echo .............. TRAN1.............
     *tran dt tstop
     
     tran 0.05u 1m
     
     
     let vds2q= v(5,6)
     let vds1q= v(6,7)
     let vgs2q= v(3,6)
     let vgs1q= v(2,7)
     let vg1=v(1)
     
     let vout=v(5)
     
     
     *fourier -popacenje
     *fourier f0 signal
     
     
     fourier 5k vout
     
     
     
     let vin_pp= max(v(1))-min(v(1))
     let vout_pp= max(v(5))-min(v(5))
     let av_abs=vout_pp/vin_pp
     
     print av_abs
   
   
   echo .............. TRAN2................
   
     tran 0.05u 1m
     
     let vgg_v= max(v(10))-min(v(10))
     let ig= max(i(vgg))-min(i(vgg))
     let rout=vgg_v/ig
     
     print rout
     
     
     
   
   
   
     
     
     
     
    
  .endc






 .end
