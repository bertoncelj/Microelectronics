Komentar, naslov, ....  //program ignorira prvo vrstico

    * Opis vezja
    * 1.crka: tip el. (r, c, l, m-mosfet, q-bipolar, v, i, ...)
    * sledi : ime el.
    * sledi : vozl.
    * sledi : parametri

    * k-kilo, m-mili, meg-mega, u-mikro,  ...
rs  4   5   r=4372
rd  2   3   r=8k

    *masa je vedno vozlisce 0
    *v_imeVira n+ n- dc=xx acmag=xx sin=(offset amp freq)
vin 1   0   dc=0    sin=(0, 1.2894, 1k)
vss 5   0   dc=-5
vdd 2   0   dc= 5

    *m_imeTran d g s b imeModela parametri
    *.model imeModela tipEl parametri(kp, vto, ...)

.model nmosTest nmos level=1 vto=1.4 kp=0.5m
m1  3   1   4   4 nmosTest w=1u l=1u

    *control zacne ukaz
.control
    destroy all

    echo #### vaja 1 ####

    
    echo ------OP1-------
        *delovna tocka
    op
    

    * print v(1) v(2) v(3) i(vin)
        * print all
    
        *tok skozi tranz. idq
    *print -i(vdd) i(vss) v(2,3)/@rd[r]
    
        *spremenljivke (vektorji)
    let idq=-i(vdd)
    let vdsq = v(3,4)
    let vgsq = v(1,4)
    let vout = v(3)
    print idq vdsq vgsq vout
    
    
    echo ------DC1------- 
        * enosmerna analiza
        * dc param start stop korak
    
    dc @rs[r] 1k 10k 10
    *plot -i(vdd)*1000 xlabel 'RS[ohm]' ylabel 'Idq[mA]'
    
    echo ------DC2-------
    
    dc vin -10 10 0.1 
    
    let id = -i(vdd)
    let vds = v(3,4)
    let vgs = v(1,4)
    let vout = v(3)
    
    *plot id vs vds xlabel 'Vds[v]' ylabel 'Id[A]'
    *plot vout xlabel 'Vin[v]' ylabel 'Vout[v]'
        * y vs x
    
    echo ------TRAN1------
        *tran dt            tstop
        *     časovni korak,konec
    tran 1u 5m
    
    let id = -i(vdd)
    let vds = v(3,4)
    let vgs = v(1,4)
    let vout = v(3)
    
    plot v(1) vout xlabel 'time' ylabel 'r:vin[t] g:vout[t]' 
    
    
        *fourier - popacenje
        *fourier f0 signal
    fourier 1k vout
    
        *racun ojacanja
    let vinPP = max(v(1))-min(v(1))
    let voutPP = max(v(3))-min(v(3))
    let avABS = voutPP/vinPP
    print avABS
    
    
    
    
    
.endc
    *vsak control potrebuje endc

.end

    *ukazi: echo, op, setplot, display, let, print, dc, destroy, plot, tran, fourier,
