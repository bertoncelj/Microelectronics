Vaja 5

    .include models.inc

    r_rc    2   4   r=1.46k
    r_re    6   0   r=1k
    r_rl    0   5   r=10k
    r_r1    3   2   r=178k
    r_r2    0   3   r=95k
    
    c_c1    1   3   c=100u
    c_c2    4   5   c=100u
    c_ce    6   0   c=100u
    
    v_vcc   2   0   dc=10
    v_vin   1   0   dc=0    sin=(0, 0.01, 5k)
    
    q1   4   3   7  T2n2222
    q2   4   7   6  T2n2222
    
    .control
    destroy all
        echo ########## Vaja 5 ##########

        
    .endc

    .end
