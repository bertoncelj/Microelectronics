 kometar, naslov...


  *opis vezja
  *1.crka     :tip el. (r,c,l,m -mostfet, q-bjt, v,i,...)
  *sledi      : ime el.
  *sledi      : vozl.
  *sledi      :parametri
  
  
  *masa: vozlisce 0
  *k-kilo, m-mili, meg - mega, u-mikro,...
  
  
  rs     4  5   r=4.4k
  rd     2  3   r=8k
  
  *v:imevira n+ n-  dc=xx acmag=xx  sin(offset, amplituda, frekvenca)
  
  vin   1  0  dc=0 sin=(0, 1.3, 1k)
  vdd   2  0  dc=5
  vss   5  0  dc=-5
  
  *m imeTranzistorja  d g  s c imeModela parametri
  * .model imeModela tipEl parametri(kp,vto, labda...)
  
  .model nmosTest nmos level=1  vto=1.4 kp=0.25m
  
  m1  3  1  4  4  nmostest  w=2u   l=1u
  
  
  

 *komentar
 *ukazi: echo, op, setplot, display, print, let ,dc, destroy, plot, tran, fourier, max, min, sqrt
 
 

  .control
     destroy all
     echo  ################Vaja 1################
     
     
     echo  .................OP1.................
     *delovna tocka
     op
     
     * print v(1), print v(2), print all, print vdd#branch,...
     
     *tok skozi tranzistor
     print -i(vdd) i(vss) v(2,3)/@rd[r]
     
     
     *spremenljivke (vektorji)
     let idq=-i(vdd)
     print idq
     
     let vdsq=v(3,4)
     let vgsq=v(1,4)
     let vout=(3)
     print idq vdsq vgsq vout
     
     
     
     
     echo ..................DC1..................
     * enosmerna analiza
     * dc parameter start stop korak
     
     dc @rs[r] 1k 10k 10
     
     plot -i(vdd) xlabel 'RS[ohm]' ylabel 'IDQ [A]'
     
     
     echo .............. DC2..............
     dc vin -10 10 0.1
     
     let id= -i(vdd)
     let vds=v(3,4)
     let vgs=v(1,4)
     let vout=v(3)
     
     * popraviti defoul scale pisemo vektor vs drugi vektor na x i y osi
     
     plot id vs vds xlabel 'vds[V]' ylabel 'id[A]'
     plot vout xlabel 'vin[V]' ylabel 'vout[V]'
     
     
      echo .............. TRAN1.............
     *tran dt tstop
     
     tran 10u 5m
     
     let id= -i(vdd)
     let vds=v(3,4)
     let vgs=v(1,4)
     let vout=v(3)
     
     plot v(1) vout xlabel 'time' ylabel 'r:vin(t), g:vout(t)'
     
     
     
     *fourier -popacenje
     *fourier f0 signal
     fourier 1k vout
     
     let vin_pp= max(v(1))-min(v(1))
     let vout_pp= max(v(3))-min(v(3))
     let av_abs=vout_pp/vin_pp
     
     print av_abs
   
  .endc






 .end
