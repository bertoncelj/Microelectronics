*test
r_rs 9 2 r=5.45k
r_rd 4 5 r=12.55k
r_r1 2 3 r=37.45k
r_r2 4 3 r=150.42k
r_si 6 7 r=500
c1  3 6 c=100u
m1 5 3 1 1 testmodel w=1u l=1u
.model testmodel pmos vto=-0.5 kp=7.5m  lambda=0
v_1 2 0  dc=9
v_2 4 0  dc=-9
v_vin 7 0 dc=0 sin=(0,2.649,5k)
c2 5 8 c=100u
rl 8 0 r=10k
v_3 1 9 dc=0
.control
destroy all
echo ...DC analiza
op
let idq=-i(v_3)
let vsd=v(1,5)
let vsg=v(1,3)
print idq vsd vsg
dc @@testmodel[kp] 7.25m 8.25m 0.1m
let idqq=-i(v_3)
plot idqq
deltaI=max(idqq)-min(idqq)
print deltaI
echo ...tran
tran 1u 1m
let vout=v(8)
let vin=v(7)
plot vout vin
echo ..fourier
fourier 5k vout 
let vin_pp=max(vin)-min(vin)
let vout_pp=max(vout)-min(vout)
let av_abs=vout_pp/vin_pp
print av_abs
.endc
.end
