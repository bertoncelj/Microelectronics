 
v_vin   1   0   dc=0    sin=(1,1,1), acmag=1
r_r1    1   2   r=1k
c_c1    2   3   c=1u
r_r2    3   0   r=2k   
c_c2    3   0   c=0.1n
 
    .control
        destroy all
        echo    ###
        *malosignalni izmenični model =>porerbuje usaj 1 acmag
        * ac tip skale st_tock  fstrat  fstop
        ac  dec 10  1   100meg
        let av=v(3)/v(1)
        let av_db=db(av)
        let av_ph=ph(av)
        plot av xlabel 'f' ylabel 'Av'
        plot av_db xlabel 'f' ylabel 'Av[db]'
        plot av_ph xlabel 'f' ylabel 'Av[ph]'
        let z1=v(1)/-i(v_vin)
        let zin=abs(z1)
        plot zin
    .endc
.end
