 Komentar,naslov,opis..
 
 
 *komentar se zacne zvezdico
 *ukazi:echo,op,seplot,desgtroy,display,print,let,plot,tran,fourier,max,min
 *opis vezja
 *elementi:
 *1.crka:tip el.(r,c,l,q,m,d,v,i,..)
 *ime elementa
 *vozlisca
 *parametri
 *koncnic:k-kilo,m-mili,M IGNORIRA VELIKE CRKE,meg-mega,u-mikro,g,t,n,p,f,
 *brez enot
  
 r_rd 2 3 r=8k
 r_rs 4 5 r=4.3k
 *v n+ n- dc= xxx sin=(offset ,ampl,ferkv) acmag=xxx
 v_vin 1 0 dc=0 sin=(0,1.5,1k)
 v_vdd 2 0 dc=5
 v_vss 5 0 dc=-5
 *mosfet
 *mime d g s b-bulk 
 m_m1 3 1 4 4 testmodel  w=2u l=1u
 *model:.model ime_modela tip_el parametri
 .model testmodel nmos vto=1.4 kp=0.25m lambda=0
  .control
  destroy all

 echo Start
 
   op
  *IDQ:vrd/rd=v(2,3)/rd
 * print  -i(v_vdd) v(2,3)/@r_rd[r]  v_vss#branch
let idq=-i(v_vdd)
let vdsq=v(3,4)
let vgsq=v(1,4)
let vout=v(3)
 print idq vdsq vgsq
 *enosmerna analiza
 echo ...........DC1......
 *dc param start stop korak
 dc @r_rs[r] 1k 10k 10
 let idq=-i(v_vdd)
let vdsq=v(3,4)
let vgsq=v(1,4)
let vout=v(3)
*plot idq xlabel 'RS[ohm]' ylabel 'IDQ [A]'

echo .....DC2...
*dc @
dc v_vin -10 10 1
let id=-i(v_vdd)
let vds=v(3,4)
let vgs=v(1,4)
let vout=v(3)
*plot id  vs vds xlabel 'vds[V]' ylabel 'i[A]'
*plot vout xlabel 'vin[V]' ylabel  'vout[v]'
echo....tran...
*tran dt stop
tran 1u 5m
 let id=-i(v_vdd)
let vds=v(3,4)
let vgs=v(1,4)
let vout=v(3)
let vin=v(1)
plot vin vout xlabel 'time' ylabel 'rvin,g:vout'
*fourier
*fourier f0 signal 
fourier 1k vout 
let vin_pp=max(vin)-min(vin)
let vout_pp=max(vout)-min(vout)
let av_abs=vout_pp/vin_pp
print av_abs
