Komentar, naslov,.....

.include models.inc


vin 1 0    dc = 0   sin=(1, 1, 5k)  acmag=1

r1 1 2     r=1k
r2 3 0     r=2k

c1 2 3 c=1u
c2 3 0 c=1n


.control
destroy all

    echo ############## AC1 ##############

    *malosignalna izmenicna analiza => potrebuje vsaj en acmag vir
    * ac tip_skale st_tock fstart fstop
    
    ac dec 100 100m 100meg
    let av      = v(3)/v(1)
    let av_db   = db(av)
    let av_ph   = ph(av)
    
    let zin     = v(1)/-i(vin)
    plot av_db xlabel 'f' ylabel 'Av[dB]'
    plot av_ph xlabel 'f' ylabel 'fi[°]'
    plot abs(zin)
    
    
    
.endc
.end
