    Komentar, naslov,..  


    * Opis vezja
    * 1. crka   : tip elementa (v pdf...r, c, t, m - mosfet,q- bjt, v, i,...=
    * sledi     : ime el.
    * sledi     : vozlisca
    * sledi     : parametri 
    
    
    
    *masa: je vedno vozlisce 0 
    * k-kilo, m-mili, meg-mega, u-mikro, n-nano, f-femto,...
    r_rs    4   5   r=4.4k
    r_rd      2   3   r=8k
    
    
    * v_imeVira n+ n- dc=xx acmag=xx sin=(offset, ampl, freq,..)
    v_vin   1   0   dc=0    sin=(0, 1.33, 1k)
    v_vdd   2   0   dc=5
    v_vss   5   0   dc=-5
    
    *m_imeTransistorja d g s b imeModela pamatri
    * .model imeModela tipElementa parametri (kp, vto, lambda,...)
    
    .model nmosTest nmos level=1 vto=1.4 kp=0.5m
    m_m1    3   1   4   4   nmosTest    w=1u    l=1u
    

    * komentar

    * ukazi: echo, op, setplot, display, print, let, dc, destroy, destroy all, plot, tran, fourier, max, min, sqrt


    .control
        destroy all
        
        
        echo ######## Vaja 1 #########
        
    
        echo --------  OP1 ------------
        * Delovna tocka
        op
        
        * print v(1) v(2) v_vin#branch i(v_vdd)
        * print all
        
        * tok skozi tranzistor IDQ
        * print -i(v_vdd) i(v_vss) v(2,3)/@r_rd[r]
        
        * spremenljivke (vektorji)
        let idq=-i(v_vdd)
        let vdsq=v(3,4)
        let vgsq=v(1,4)
        let vout=v(3)
        print idq vdsq vgsq vout
        
        
        
        echo --------  DC1 ------------
        * Enosmerna analiza
        * dc parameter start stop korak
        dc @r_rs[r] 1k 10k 10
        
        *plot -i(v_vdd) xlabel 'RS[ohm]' ylabel 'IDQ [A]'
        
        
        echo --------  DC2 ------------
        dc v_vin -10 10 0.1
        
        let id=-i(v_vdd)
        let vds=v(3,4)
        let vgs=v(1,4)
        let vout=v(3)
     
        
        *plot id vs vds xlabel 'vds[V]' ylabel 'id[A]'
        *plot vout xlabel 'vin[V]' ylabel 'vout[V]'
        
        
        
        echo --------  TRAN1 ------------
        * tran dt tstop -> dt-casovni korak, da je pokritost periode 100, 1000 tock, tstop-cas analize
        tran 10u 5m 
        
        let id=-i(v_vdd)
        let vds=v(3,4)
        let vgs=v(1,4)
        let vout=v(3)
        
        plot v(1) vout xlabel 'time' ylabel 'r:vin(t), g:vout(t)'
        
        
        * fourier - popacenje
        * fourier f0 signal
        fourier 1k vout
        
        
        let v_in_pp=max(v(1))-min(v(1))
        let v_out_pp=max(v(3))-min(v(3))        
        let av_abs=v_out_pp/v_in_pp
        
        print av_abs
        
        
    .endc

    .end
