Moje prvo vezje
v1 1 0 dc=5
r1 1 2 r=40.4864k
r2 3 2 r=31.63k
r3 3 4 r=54.4k
v2 4 0 dc=-5
v3 7 8 dc=0
rs 4 5 r=5k
rd 8 1 r=5k
c1 3 9 c=1u
v_vin 9 0 dc=0 sin=(0,0,0)
vx 11 0 dc=0 sin=(0,0.201,5k)
c4 7 10 c=100u
v4 10 11 dc=0
c2 2 0 c=100u
c3 5 0 c=100u
m1 7 2 6 6  testmodel 
m2 6 3 5 5 testmodel 
.model testmodel nmos vto=0.8 kp=1m  lambda=0
.control
op
echo ...op
let vdsq2=v(7)-v(6)
let vdsq1=v(6)-v(5)
let idq=-i(v3)
let vgs2=v(2)-v(6)
let vgs1=v(3)-v(5)
let Vg1=v(3)
print Vg1 vdsq2 vdsq1 idq vgs2 vgs1
echo ...tran
tran 1u 1m
let ix=i(vx)
ixpp=max(ix)-min(ix)
vxpp=max(v(11))-min(v(11))
rout=vxpp/ixpp
print rout
.endc
.end
