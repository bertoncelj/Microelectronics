3.Lab Vaja: MOSFET  kaskodni ojačevalnik
*Tf je funkcija ki iz vefje izpljuune vn kondeznatorje
*ampak se jo ne rabi pri linearni elektroniki
 
   	*upornosti
    r_r1    1   2   r=40.5k
    r_r2    2   3   r=31.6k
    r_r3    3   4   r=54.4k
    
    r_rs    5   4   r=5k
    r_rd    1   8   r=5k
    
    *kapacitiovnosti
    c_c1    10    3    c=100u
    c_c2    2    0     c=100u
    c_c3    5    0     c=100u
    
    *napajalniki
    v_plus    1   0   dc=5     
    v_minus   4   0   dc=-5
    v_vg_in   9   0   dc=0 sin(0, 201m, 5k) 
    *amplitudna vrednost sinusa se probava, da gledas vrednost THC procent  napake!
    
    *dodamo merilni napajalnik
    vmer 9 10 dc = 0
    
    * m_imeTran d g s b (drain, gate, source, base) imeModela parametri
   .model nmos_model nmos level=1 vto=0.8 kp=1m
    m_m1    6   3   5   5   nmos_model    w=1u    l=1u
    m_m2    8   2   6   6   nmos_model    w=1u    l=1u
   
    .control
        destroy all
        
        echo _______________VAJA 2______________
        echo 
        
        *naredi DC analizo
        op

        *nastavimo vektorje ki jih iscemo
        let idq= v(5,4)/@r_rs[r]
        let vdsq1 = v(8,6)
        let vdsq2 = v(6,5)
        let vgsq1 = v(3,5)
        let vgsq2 = v(2,6)
        let vg1   = v(2)
        
        *izise vse nastavljene vektorje ki jih gledamo
        print idq vdsq1 vdsq2 vgsq1 vgsq2 vg1
        
        echo _______________VAJA 3______________
        echo

        tran 1u 2m
        
        *dolocimo vektorje 
        let vin  = v(3)
        let vout = v(8)
        
        *izrise graf
        * plot vin vout v(6) xlabel 'time' ylabel 'vg1, vd2, vs1'
        *plot vin vout xlabel 'time [s]' ylabel 'r:vin(t), g:vout(t)'
         
        fourier 5k vout
        
        let vin_PP = max(vin)-min(vin)
    	let vout_PP = max(vout)-min(vout)
        
        let av = vout_PP/vin_PP
        echo ___________HERE________________
        let rin = vin_PP/(max(i(vmer))-min(i(vmer)))
        echo ___________HERE_______________
        let rout = vout_pp/((max(v(1,8))-min(v(1,8)))/@r_rd[r])
        echo ___________HERE_______________
        
        print av rin rout
         
         echo _______________VAJA 4______________
        echo
         *Casovna analiza
         
         
    .endc
    
.end
