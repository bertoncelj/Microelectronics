vaja 3

*.include models.inc

	vin 	1 0 dc=0 sin=(0, 0.5166, 5k)
	vp 		5 0 dc=5
	vn 		4 0 dc=-5
	vtest	8 5 dc=0
	r1 		3 5 r=242k
	r2 		3 4 r=395k
	re		4 6 r=10k
	*rl		7 0 r=2.000k
	rsrc	1 2 r=10.000k
	rl		7 0 r=20.000k
	c1 		2 3 c=100u
	c2 		6 7 c=100u
	
	
	
	q (8 3 6 )   BC238B 
	
.MODEL BC238B NPN IS=1.8E-14 ISE=5.0E-14 NF=.9955 NE=1.46 BF=400 BR=35.5
+ IKF=.14 IKR=.03 ISC=1.72E-13 NC=1.27 NR=1.005 RB=.56 RE=.6 RC=.25 VAF=80
+ VAR=12.5 CJE=13E-12 TF=.64E-9 CJC=4E-12 TR=50.72E-9 VJC=.54 MJC=.33

	



.control
	destroy all


    op
	let icq=-i(vtest) 
	let vceq=v(8,6)
	let vbeq=v(3,6)
	print icq vceq vbeq
	
	tran 1u 5m
	let vout=v(7)
	let vin=v(1)
	let vin_pp=max(vin)-min(vin)
	let vout_pp=max(vout)-min(vout)
	let av=vout_pp/vin_pp
    plot vin vout
	print  av
	
	fourier 5k vout
	let iout=v(7)/@rl[r]
	let iin=v(1,2)/@rsrc[r]
	let iin_pp=max(iin)-min(iin)
	let iout_pp=max(iout)-min(iout)
	let ai=iout_pp/iin_pp
	
	print ai
	
.endc
.end
