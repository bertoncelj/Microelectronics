2. Laboratorijska vaja

*OPIS VEZJA

	vin 7 0 dc=0 sin=(0, 0.0140, 5k)
	vp 1 0 dc=9
	vn 0 3 dc=9

	rsi 7 8 r=500
	r1 1 2 r=37.5k
	r2 2 3 r=150.8k
	rs 1 5 r=5432
	rd 4 3 r=12551.5
	rl 6 0 r=10k

	c1 8 2 c=100u
	c2 4 6 c=100u
	cs 5 0 c=100u

	m1 4 2 5 5 testmodela w=15u l=1u 
	.model testmodela pmos vto=-0.5 kp=0.55m lambda=0

.control
destroy all
	echo ############DRUGAVAJA#######

	echo -----------DelovnaTocka--------------

	op
		let idq=v(1,5)/@rs[r]
		let vsdq=v(5,4)
		let vsgq=v(5,2)
		print idq vsdq vsgq
		
	echo ------------tran1----------

	tran 0.5u 5m
	
	let id=v(1,5)/@rs[r]
	let vsd=v(5,4)
	let vsg=v(5,2)
	let vout=v(6)
	let vin=v(7)
	let vss=v(5)
	let vgg=v(2)
	let vdd=v(4)

	fourier 5k vout
	plot vss vgg vdd xlabel 'time' ylabel 'vs, vg, vd'

	let vin_pp=max(vin)-min(vin)
	let vout_pp=max(vout)-min(vout)
	let av=vout_pp/vin_pp

	vss_pp=max(vss)-min(vss)
	vgg_pp=max(vgg)-min(vgg)
	vdd_pp=max(vdd)-min(vdd)

	print av vss_pp vgg_pp vdd_pp
.endc
.end
	
