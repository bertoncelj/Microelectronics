 Komentar, naslov, opis vezja, ...
 .include models.inc
 * Komentar se začne z zvezdico in obsega celo vrstico
 
 * Opis vezja
 * Elementi:
 * 1. crka: Tip elementa (r, c, l, q, m, d, v, i, ...)
 * sledi: ime elementa
 * sledi: vozlisca
 * sledi: parametri
 * Koncnice potenc 10: k-kilo, m-mili, meg-mega, u-mikro, g-giga, t-tera, n-nano
 * Brez enot
 
*-----------------------------------------------------------------------------------------------------
	
	r1		3	4	r=242k
	r2		3	6	r=395k
	re		5	6	r=10k
	rl		7	0	r=20k
	rsrc	1	2	r=10k
	
*-----------------------------------------------------------------------------------------------------
	
	c1	2	3	c=100u
	c2	5	7	c=100u
		
*-----------------------------------------------------------------------------------------------------
 * v_ime        n+  n-  dc=xxx 	sin=(offset, amplituda, frekvenca)   acmag=xxx
 
	vsrc 		1	0 	dc=0 	sin=(0, 0.2010767, 5k)
	vp 			4 	0 	dc=5
	vn 			6 	0 	dc=-5

*-----------------------------------------------------------------------------------------------------

* Mosfet
 * m_ime        drain   gate   source   bulk    ime_modela  parametri
	*m1			4		3	   5        5       BC238B   	
	
* Bipolarni
 * q_ime        colector    base    emitor      ime_modela
    q1          4           3       5           BC238B
*-----------------------------------------------------------------------------------------------------	

* model: .model 	ime_modela 	tip_elementa 	parametri (kp parameter je v ucbeniku kp')	
		 .model 	testmodel   nmos      		vto=0.8 kp=0.5m lambda=0.0001
		 
*-----------------------------------------------------------------------------------------------------

* Kontrol blok, notri so ukazi
* Ukazi: echo (izpiše tekst v okno simulatorja)
*        cd (zamenja mapo)
*        op (analiza delovne tocke)
*        setplot
*        destroy (all ali posamezno)
*        display (pokaze kaj je SPICE izracunal v zadnji analizi)
*        i(ime vira) (dostop do toka skozi vir)
*        let (to je za delat s spremenljivkami)
*        dc (dc analiza)
*        plot ()
*        tf  out vir
		 
*-----------------------------------------------------------------------------------------------------

.control																		
    destroy all																	
																				
	echo ###########################START############################
    
	echo --------------------------__OP1__---------------------------
    
	op
			
			let beta = 150
			let icq = v(5,6)/@re[r]*((beta-1)/beta)
			let vceq = v(4,5)
			let vbeq = v(3,5)
			
			print icq vceq vbeq
	
	echo --------------------------_TRAN1_---------------------------
		
		tran 1u 5m
			
			let icq = v(3,4)/@r1[r]
			let vceq = v(4,5)
			let vbeq = v(3,5)
			
			let vout=v(7)
			let vsrc=v(1)
			let vp=v(4)
			let vn=v(8)
			
			fourier 5k vout
			*plot vin vout xlabel 'cas' ylabel 'Vin[V] - red	  Vout[V] - green'
			
			let vsrc_pp=max(vsrc)-min(vsrc)
			let vout_pp=max(vout)-min(vout)
			let av=-vout_pp/vsrc_pp
			
			print av
			
			*let isrc_pp = max(i(vsrc))-min(i(vsrc))
			*let vx_pp = max(v(2,8))-min(v(2,8))
			*let rin = vx_pp/iin_pp
			
			*print rin
			
			*let iout_pp = max(i(vx))-min(i(vx))
			*let rout = vout_pp/iout_pp
			
			*print rout
			
	.endc

.end

*-----------------------------------------------------------------------------------------------------


* Dostop do vaj od doma: lisa.fe.uni-lj.si/vaje    Uporabnik: vaje Geslo: vajenec
