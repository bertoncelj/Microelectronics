Komentar, naslov, opis, ...

* komentarji z zvezdico


* opis vezja
* elementi:
*   1. crka: rip el. (rm cm l, q, m, d v, i, ...)
*   sledi: ime el.
*   sledi: vozlišča

* koncnice potenc 10: f, p, n, u, m, k, meg, g, t
* brez enot!

r_rd 2 3 r=8k
r_rs 4 5 r=4.37k

* v_ime n+ n- dc=xxx sin=(offset, ampl, frekv) acmag=xxx
v_vin 1 0 dc=0 sin=(0, 1, 1k)
v_vdd 2 0 dc=5
v_vss 5 0 dc=-5


* mosfet
* m_ime drain gate source bulk ime_modela parametri
m_m1 3 1 4 4 testmodel w=2u l=1u

* model: .model ime_modela tip_el parametri
* Kn = 1/2 * kn' W/L <-- spice opus uporablja kn' oz. kp
* če navodilo 0.25mAV^-2, sami ustrezno zložimo parametre
* pod model pišemo lastnosti tehnologije, pod m pa posameznega tranzistorja
.model testmodel nmos vto=1.4 kp=0.25m lambda=0


* ampermeter v spicu: avt. racuna tok. dolocimo v_m1 dc=0 --> dobimo tok

* IDQ = Kn(VGSQ - VTN)^2 --> VGSQ = ...
* -VinDC (je 0) + VGSQ + IDQ*RS + VSS = 0 --> Rs = ...
* IDQ = (VDD - VOUT) / RD --> RD = 8kOhm
* IDQ*RD + IDSQ + IDQ*RS + VSS - VDD = 0 --> VDSQ = ... > VDS,sat = UGSQ - VTN (sicer lin.)


* konrol block - ukazi
* ukazi: echo, op, setplot, destroy, display, print, plot, ttran, fourier, max, min, let, dc

.control
    destroy all

    echo ######## START ########

    echo --------- OP1 ---------
    op

    * IDQ: vRD/RD = v(1,2)/rd
    *print v(2,3)/@r_rd[r]
    *print -i(v_vdd)
    *print v_vss#branch

    let idq = -i(v_vdd)
    let vdsq = v(3,4)
    let vgsq = v(1,4)
    let vout = v(3)
    
    print idq vdsq vgsq vout
    

    *enosmerna analiza
    echo --------- DC1 ---------
    * dc param start stop korak
    dc @r_rs[r] 1k 10k 10
    
    let idq = -i(v_vdd)
    let vdsq = v(3,4)
    let vgsq = v(1,4)
    let vout = v(3)
    
    *plot idq xlabel 'RS [ohm]' ylabel 'IDQ [A]'
    
    echo --------- DC2 ---------
    *DC @v_vin[dc] -10 10 1
    dc v_vin -10 10 0.1
    
    let id = -i(v_vdd)
    let vds = v(3,4)
    let vgs = v(1,4)
    let vout = v(3)
    
    *plot id xlabel 'vin[V]' ylabel 'id[A]'
    *plot id vs vds xlabel 'vds[V]' ylabel 'id[A]'
    *plot vout vs sweep xlabel 'v[V]' ylabel 'vout[V]'
    
    echo -------- TRAN1 --------
    * tran dt tstop
    tran 1u 5m
    
    let id = -i(v_vdd)
    let vds = v(3,4)
    let vgs = v(1,4)
    let vout = v(3)
    let vin = v(1)
    
    *plot vin vout xlabel 'time' ylabel 'r:vin, g:vout'
    
    
    * fourier - analiza popačenja
    * fourier f0 signal
    fourier 1k vout
    
    let vin_pp=max(vin)-min(vin)
    let vout_pp=max(vout)-min(vout)
    let av_abs=vout_pp/vin_pp
    print av_abs
    
.endc

.end
