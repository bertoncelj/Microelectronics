Vaja 3 kaskodna vezava nMos


vp 		5 	0 	dc = 5
vn 		7 	0 	dc = -5
vin 	8 	0 	dc = 0	sin=(0, 0, 5k) 
vtest   10  0   dc=0 sin=(0,1,5k)
r1 	3 	5	r=40.5k
r2 	1 	3 	r=31.6k
r3 	7 	1 	r=54.4k
rs 	6 	7 	r=5k
rd 	5 	4 	r=5k

c1	 8	 1 	c=100u
c2	 3	 0 	c=100u
c3	 6	 0 	c=100u
c4   4  10  c=100u
	*m_imeTran d g s b imeModela parametri
	*.model imeModela tipEl parametri(kp, vto, ...)

.model modeln nmos kp=0.5m vto=0.8 lambda=0.1m

m1 2 1 6 6 modeln w=2u l=1u
m2 4 3 2 2 modeln w=2u l=1u	
	

.control
destroy all
    

    
    echo ---------OP1---
	op
	let idq = v(5,4)/5000
	let vdsq1 = v(2,6)
	let vdsq2 = v(4,2)
	let vgsq1 = v(1,6)
	let vgsq2 = v(3,2)
	let vg1	  = v(1)
	
	print idq vdsq1 vdsq2 vgsq1 vgsq2 vg1 
	
	
	
	
	
	
	echo ---------tran--
	
	tran 1u 5m
    
    let vin=v(8)
    let vout=v(10)
    
    
    
    
    let vin_pp=max(vin)-min(vin)
    let vout_pp=max(vout) - min (vout)
    let av_abs=vout_pp/vin_pp
    let rout = vout_pp/((max(v(4,5))-min(v(4,5)))/5000)
    print  rout
	
	
	
    
.endc
.end
