 4. Laboratorijska vaja (Komentar,naslov,....)

    .include models.inc
 
    *Ukazi: echo, op(delona tocka), setplot, display, print, let, dc, destroy, plot, tran, fourier, max, min
    *-------opis vezja------------------
	
	
    r_re    6   0   r=1k
	r_r1    3   2   r=178k
	r_r2    2   0   r=95k
	r_rl    7   0   r=10k
    r_rc    3   4   r=1.46k
    

	v_vin   1   0   dc=0    sin=(0, 0.20, 5k), acmag=1
    v_vcc   3   0   dc=10
    v_vmer1 4   441  dc=0
    v_vmer2 4   442  dc=0
	
	q_q1   441   2   5   T2N2222
	q_q2   442   5   6   T2N2222
	
	
	C1     1	2	c=100u	
	C2     4	7	c=100u	
	ce     6    0   c=100u
	
	*------------Simulacija-----------------
    
    .control
        destroy all
    
        echo ######### Vaja 5 #########
        
        
        echo --------- op1 ---------
		
		*delovna tocka
		op
		
        let vceq1=v(4,5)
        let vceq2=v(4,6)
		let icq1=i(v_vmer1)
		let icq2=i(v_vmer2)
		
		
        print vceq1 vceq2 icq1 icq2
        
        echo --------- TRAN1 ---------
        
		* tran dt tstop --- casovna analiza (dt-CASOVNI korak, )
		

        
        
    .endc

    .end
 
