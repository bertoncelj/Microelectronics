Komentar, naslov,..... kar napišeš v prvi vrstici spice ignorira


*OpisVezja:
*1.crka: tip elementa (r, c, l, m - mos tranzistor, q- bipolarc, v - napet vir, i tok vir,....)
*      : ime elementa
*      : vozlisca
*      : parametri

* k- kilo, m - mili, meg - mega, u- mikro.....

rs  4   5   r=500k
rd  2   3   r=5k


*v_imeVira n+ n- parametri: dc= neki, acmag= neki sin=(neki) vedno najprej pozitivno

vin 1   0   dc=0
vdd 2   0   dc=5
vss 5   0   dc=-5

*m_imeTran d g s b (vrstni red je pomemben) ime modela parametri
*.model imeModela tipElementa parametri (kp, vto, lambda,....)

.model nmosTest nmos level=1 vto=1.4 kp=0.5m
m1  3   1   4   4   nmosTest    w=1u    l=1u


*komentar 
*ukaz: echo, 

.control
    echo ##################### VAJA ######## 
    
    echo ------------ OP1 -----------

    echo ------------ DC1 -----------
    
    
.endc


.end
