 


.include models.inc

vp 4 0 dc = 5
vn 5 0 dc = -5
vin 1 0 dc = 0 sin=(0, 0.1, 5k)


r1  2 4    r=242k
r2  2 5    r=395k
re  3 5    r=10k
rsrc 1 8   r=10k
rl 6 0 r=2k

c1 8 2 c=100u
c2 3 6 c=100u



q1 4 2 3 BC238B  
	

.control
destroy all
    echo ----------------------------------------------  
    
    tran 0.05 1m
    
    
   
     let Avo= max(v(6))-min(v(6))
     let Avi= max(v(8))-min(v(8))
     
     let Aio= (max(v(6))-min(v(6)))/20k
     let Aii=  max(i(vin))-min(i(vin))
     
     let Av= Avo/Avi
     let Ai= Aio/Aii
   
   
   
   print Av Ai
    
    
     
    
.endc
.end
