Naloga 2

    *DC analiza
    *vhodni
    r_r1    1   2   r= 37.4k
    r_r2    2   5   r= 151.5k
    
    
    r_rs    1   3   r= 5.4k
    r_rd    4   5   r= 12.6k
    
    *napajalniki
    v_vgate      2   0   dc=  5.436      
    v_vplus      1   0   dc=  9
    v_vminus     5   0   dc= -9
    
  * m_imeTran d g s b (drain, gate, source, base) imeModela parametri
    * .model imeModela  tipElementa parametri(kp, vto, lambda,..)
    
    .model pmosTest pmos level=1 vto=-0.5 kp=0.5m
    m_ml    4   2   3   3   pmosTest    w=15u    l=1u
    
    .control
        
        echo /************** VAJA 2 ******************/
        *pobrisemo vse spremeljivke, prosti polnilnik
        destroy all
        
        *delovna tocka op -> poisce delovno tocko
        op
        
        * tok skozi tranzistor
        print -i(v_vplus) i(v_vminus)    v(4,5)/@r_rd[r]
        
        *dolocimo numericno stevilke
        let idq  = v(1,3)/@r_rs[r]
        let vsdq = v(3,4)
        let vsgq = v(3,2)
        let vout = v(4)
        
        *izpis stevilk
        print idq vsdq vsgq vout
        
        
        
        
        
        
      .endc
 .end

