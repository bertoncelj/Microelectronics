 
.include models.inc



vcc 2 0 dc = 10
vin 1 0 dc = 0	sin=(0, 0.01, 5k)

r1 3 2 r=178k
r2 3 0 r=95k
re 6 0 r=1k
rl 5 0 r=10k
rc 2 4 r=1.46k

c1 1 3 c=100u
c2 4 5 c=100u
ce 6 0 c=100u


q1 4 3 7 T2n2222
q2 4 7 6 T2n2222

*cbe ime modela


.control
destroy all
    echo #### Vaja 5 ####

    
    echo ------OP1-------
	op
	let irc = v(2,4)/1460
	let icq1 = irc/101
	let icq2 =100*icq1 
	let vceq1 = v(4,7)
	let vceq2 = v(4,6)

	print icq1 vceq1 vceq2 icq2  
	
	
	
	echo ------TRAN1------
	
    tran 1u 5m
    let vin =v(1)
    let vout=v(5)
    let vinPP = max(v(1))-min(v(1))
    let voutPP = max(v(5))-min(v(5))
    let av = voutPP/vinPP
    print av
    
    let iin1 = max(i(vin))-min(i(vin))
    let iout1 = max(v(5)/10000)-min(v(5)/10000)
    let ai = iout1/iin1

print ai
.endc
 
.end
