asdf
 
	.include models.inc
	r1		3	4	r=242k
	r2		3	5	r=395k
	re		5	6	r=10k
	*rl		7	0	r=20k
	vx     7   0   dc=0 sin=(0,1,5k)
	rsrc	1	2	r=10k
	
	c1	2	3	c=100u
	c2	6	7	c=100u
 
	vsrc 		1	0 	dc=0
	vp 			4 	0 	dc=5
	vn 			5 	0 	dc=-5
    
    q 4 3 6 BC238B
	
*q_q1 c b e model
	
.control																		
    destroy all																	
																				
	echo ###########################START############################
    
	echo --------------------------__OP1__---------------------------
    
	op
			
			let B = 150
			let icq = v(5,6)/@re[r] *(B-1)/B
			let vceq = v(4,6)
			let vbeq = v(3,6)
			
			print icq vceq vbeq
	
	echo --------------------------_TRAN1_---------------------------
		
		tran 1u 5m
			
			let B = 150
			let icq = v(5,6)/@re[r] *(B-1)/B
			
			*fourier 5k vout
			
			*plot vin vout xlabel 'cas' ylabel 'Vin[V] - red	  Vout[V] - green'
			
			let iout_pp = max(i(vx))-min(i(vx))
			let rout = 2/iout_pp
			
			print rout
			
	.endc

.end

