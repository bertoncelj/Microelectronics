Komentar, naslov,.....

.include models.inc

vp 3 0 dc = 5
vn 4 0 dc = -5
vin 6 0 dc = 0 sin=(0, 0.1, 5k)

r1 3 1      r=242k
r2 1 4      r=395k
rsrc 6 5    r=10k
re 2 4      r=10k
rl 7 0      r=2k

c1 5 1 c=100u
c2 2 7 c=100u


q1 3 1 2 BC238B  
	

.control
destroy all
    echo ############## OP ##############
    
    op
    let ieq  = v(2,4)/@re[r] 
    let vceq = v(3,2)
    let vbeq = v(1,2)
    let icq  = i(vp)-v(3,1)/@r1[r]
    
    print ieq vceq vbeq icq
 
    echo ############## tran1 ############### 

    tran 1u 5m
    fourier 5k v(7)
    
    
    let vinPP = max(v(6))-min(v(6))
    let voutPP = max(v(7))-min(v(7))
    let avmin = voutPP/vinPP
    
    let iout = v(7)/@rl[r]
    let iinPP = max(i(vin))-min(i(vin))
    let ioutPP = max(iout)-min(iout)
    let ai1 = ioutPP/iinPP
    
    print avmin ai1
    
    echo ############## tran2 ###############     
    let @rl[r] = 20k
    tran 1u 5m
    
    let vinPP = max(v(6))-min(v(6))
    let voutPP = max(v(7))-min(v(7))
    let avmax = voutPP/vinPP
    
    let avr = tran1.avmin/avmax
    print avr avmax
    
    let iout = v(7)/@rl[r]
    let iinPP = max(i(vin))-min(i(vin))
    let ioutPP = max(iout)-min(iout)
    let ai2 = ioutPP/iinPP
    print ai2
    
.endc
.end
