 Komentar,naslov,... prvo vrstico Spice ignorira
 
 *kar se začne z zvezdico je komentar
 * kar se začne s piko (.) je ukaz
 * ukazi: echo,op(enosmerna analiza),setplot
 *(zbirka rezultatov),print,let,dc,plot,tran,fourier,
 *max(),min(),sqrt()
 
 *opis vezja
 *1.črka    : je tip elementa (r,c,l,m(mos tranzistor),q(bipolarni *tranzistor),v,i,...)
 *sledi     : ime el.
 *sledi     : vozlišča
 *sledi     :parametri
 
 *masa je vedno vozlišče 0
 *imena vseh ostalih vozlišč niso pomembna
 *k-kilo,m-mili,meg-mega,u-mikro,...
 r_rs   4   5   r=4.38k
 r_rd   2   3   r=8k
 
 *v_imeVira n+ n-   dc=xx   acmag=xx    sin=(offset,amplituda,frekvenca)
 v_vin  1   0   dc=0    sin(0,1.33,1k)
 v_vdd  2   0   dc=5
 v_vss  5   0   dc=-5
 
 *m_ime tranzistorja    d   g   s   b   imeModela   parametri
 *.model imeModela  tipElementa parametri(kp,vto,lambda,...)
 
 .model nmosTest    nmos    level=1 vto=1.4 kp=0.25m
 
 m_m1   3   1   4   4   nmosTest    w=2u    l=1u
 
 .control
    
    destroy all
    
    echo ##################### Vaja 1 ############################
    
    
    echo ---------------------- OP1 -----------------------------
    *Delovna točka
    op
    
   * print v(1) v(2) v_vin#branch i(v_vdd)
    *print all
    
    *tok skozi tranzistor IDQ
    *print -i(v_vdd) i(v_vss) v(2,3)/@r_rd[r]
    
    *spremenljivke (vektorji)
    let IDQ=-i(v_vdd)
    let VDSQ=v(3,4)
    let VGSQ=v(1,4)
    let vout=v(3)
    print idq vdsq vgsq vout
     echo ---------------------- DC1 -----------------------------
     
     *enosmerna analiza
     *dc    parameter   start   stop    korak
     
     dc     @r_rs[r]    1k      10k     10
     
     *plot -i(v_vdd) xlabel 'RS[ohm]' ylabel 'IDQ[A]'
    echo ---------------------- DC2 -----------------------------
    dc v_vin -10 10 0.1
    
    let id=-i(v_vdd)
    let vds=v(3,4)
    let vgs=v(1,4)
    let vout=v(3)
    
    *plot id vs vds xlabel 'vds[V]' ylabel 'id[A]'
    *plot vout xlabel 'vin[V]' ylabel 'vout[V]'
    
     echo ---------------------- TRAN1 -----------------------------
     
    
    
    
    *tran dt tstop
    
     
    
    
    tran 10u 5m
    
    let id=-i(v_vdd)
    let vds=v(3,4)
    let vgs=v(1,4)
    let vout=v(3)
    let vin=v(1)
    
    plot vin vout xlabel 'time' ylabel 'vin(t),vout(t)'
    
    *fourier -popačenje (mora biti znootraj transientne analize
    *fourier f0 signal
    fourier 1k vout
    
    let vin_pp=max(v(1))-min(v(1))
    let vout_pp=max(v(3))-min(v(3))
    let av_abs=vout_pp/vin_pp
    print av_abs
     
 .endc
 
 
 .end
