Emitorski sledilnik
.include models.inc

vin 1 0 dc = 0
vp 6 0 dc = 5
vn  4 0 dc = -5
vout 7 0 dc = 0 sin(0 1 5k)

r1 6 3 r=242k
r2 3 4 r=395k
re 4 5 r=10k

rsrc 1 2 r=10k

q1 6 3 5 BC238B

c1 2 3 c=100u
c2 5 7 c=100u

.control

echo ##### izhodna upornost########
echo ---------- tran -------

tran 1u 2m

let ix = max(i(vout)) - min(i(vout))
let vx = max(v(7)) - min(v(7))
let rout = vx/ix

print rout



.endc
.end
