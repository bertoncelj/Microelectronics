.include models.inc

vin 1 0 dc = 0	sin=(0, 0, 5k)
vp 6 0 dc = 5
vn 4 0 dc = -5
vx 7 0 dc = 0   sin=(0, 0.2, 5k)

r1 6 3 r=242k
r2 3 4 r=395k
re 4 5 r=10k
rsrc 1 2 r=10k

c1 2 3 c=100u
c2 5 7 c=100u

q1 6 3 5 BC238B

*cbe ime modela


.control
destroy all
	
	
	echo ------TRAN1------
	
    tran 1u 5m
    
    let vxPP = max(v(7))-min(v(7))
    let ixPP = max(i(vx))-min(i(vx))
	let rout = vxPP/ixPP
	
	print rout
	
.endc
.end
