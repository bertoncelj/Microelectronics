 Primer za 5to vajo

 
    *-------opis vezja------------------
    

	
	vin    1   0   dc=0 sin=(1,1,1k), acmag=1
	r1     1   2   r=1k
	c1     2   3   c=1u
	r2     3   0   r=2k
	c2     3   0   c=0.1n
	
	

	
	*------------Simulacija-----------------
    
    .control
    destroy all
		
            echo ######### ac analiza ###########
            * Malosignalna izmenicna analiza
            *vzbujanje za ac analizo je acmag!!
            * ac tip_skale st_tock fstart fstop
            
            ac  dec 10  1   100meg
            
            let av=v(3)/v(1)
            let av_db=db(av)
            let av_ph=ph(av)
            
            plot av_db xlabel 'f' ylabel 'Av[dB]'
            plot av_ph xlabel 'f' ylabel 'faza'
            
		
    .endc

    .end
 
