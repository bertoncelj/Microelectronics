Komentar, naslov....(SPICE ignorira)
    
    *OPIS VEZJA
    *prva črka tip rl. (r, c, l, m-mosfet, v, i ...)
    *sledi ime elementa
    *sledi vozlišča
    *sledi parametri
    
    *masa je vedno vzlisce 0
    *k-kilo, m-mili, meg-mega, u-mikro
    r_r1    3   4   r=45.6k
    r_r2    3   2   r=35.625k
    r_r3    2   5   r=61.275k
    r_rs    5   6   r=5k
    r_rd    4   7   r=5k
    
    c_c1    1   2   c=100u
    c_c2    3   0   c=100u
    c_c3    6   0   c=100u
    c_c5    7   10  c=100u
    
    *v_imevira  n+   n- dc=xx   acmag=xx    sin=(off, amp, freq)
    v_vin   1   0   dc=0   sin=(0, 0, 5k)  
    v_vp    4   0   dc=5
    v_vm    5   0   dc=-5
    v_out   10  0   dc=0    sin(0,0.1,5k)
    
    *m_imeTranz d   g   s   b   incModela parametri
    *. model imeModela tipEl parametri (kp, vto, lambda...)
    .model  nmosTest    nmos    level=1    vto=0.8  kp=0.5m

    m_m1    7   3   8   8   nmosTest    w=2u    l=1u
    m_m2    8   2   6   6   nmosTest    w=2u    l=1u
    
    *komentar
    *ukazi: echo, op, setplot(zbirka rezultatov), display, print, let,dc, destroy all, plot. tran, fourier, max, min, sqrt
     
     .control
        destroy all
        echo ######## Vaja3 ######
        echo ---------OP1---------
        *delovna tocka ukaz op
        op
        *spremenljivka (vektor)
        let idq=v(4,7)/@r_rd
        let vdsq1=v(7,8)
        let vdsq2=v(8,6)
        let vgsq1=v(3,8)
        let vgsq2=v(2,6)
        let vg1=v(2)
        let iout=i(v_vout)
        print idq, vdsq1, vdsq2, vgsq1, vgsq2, vg1 ,
        echo -------TRAN1-------
        tran 1u 5m
       * fourier 5k v(7)
        echo -------TRAN2-------
        *let vin_pp = max(v(1))-min(v(1))
        let vout_pp = max(v(7))-min(v(7))
        let iout_pp=max(i(v_out))-min(i(v_out))
        *let Av=vout_pp/vin_pp
        let rout=vout_pp/iout_pp
        print rout
        
    .endc
    
    .end

